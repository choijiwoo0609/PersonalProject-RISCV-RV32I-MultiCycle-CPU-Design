`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:50];

    initial begin
        //$readmemh("code.mem", rom);

        //rom[x]=32'b  funct7_ rs2 _ rs1 _ f3 _ rd _ op       // R-Type                  rd   |    r1    |   r2  
        rom[0] =  32'b0000000_00001_00010_000_00011_0110011;  // add  x3, x2, x1  =>     23   |    12    |   11             
        rom[1] =  32'b0100000_00001_00010_000_00100_0110011;  // sub  x4, x2, x1  =>      1   |    12    |   11        
        rom[2] =  32'b0000000_10010_00010_001_00101_0110011;  // sll  x5, x2, x18 => 1100..00 |    12    |   28    -> signed로 볼 경우 : 3221225472 / unsigned로 볼 경우 : -1073741824
        rom[3] =  32'b0000000_00001_00010_101_00110_0110011;  // srl  x6 x2, x1   =>      0   |    12    |   11        
        rom[4] =  32'b0100000_00001_00010_101_00111_0110011;  // sra  x7 x2, x1   =>      0   |    12    |   11        
        rom[5] =  32'b0000000_00010_00101_010_01000_0110011;  // slt  x8 x5, x2   =>      1   | (-107...)|   12    -> signed 이므로 1이 출력됨      
        rom[6] =  32'b0000000_00010_00101_011_01001_0110011;  // sltu x9 x5, x2   =>      0   | (3221...)|   12    -> unsigned 이므로 0이 출력됨.    
        rom[7] =  32'b0000000_00010_00001_100_01010_0110011;  // xor  x10 x1, x2  =>  7(0111) | 11(1011) | 12(1100)        
        rom[8] =  32'b0000000_00010_00001_110_01011_0110011;  // or   x11 x1, x2  => 15(1111) | 11(1011) | 12(1100)        
        rom[9] =  32'b0000000_00010_00001_111_01100_0110011;  // and  x12 x1, x2  =>  8(1000) | 11(1011) | 12(1100)        
  
        //rom[x]=32'b    imm12    _ rs1 _ f3_ rd  _ op       // I-TYPE (12-bit immediate)      rd   |   r1     |   imm      
        rom[10] = 32'b000000000001_00010_000_00110_0010011;  // addi x6, x2, 1           =>    13   |   12     |     1              
        rom[11] = 32'b000000000001_00101_010_00111_0010011;  // slti x7, x5, 1           =>     1   | (-107...)|     1        -> signed 이므로 1이 출력됨    
        rom[12] = 32'b000000000001_00101_011_01000_0010011;  // sltiu x8, x5, 1          =>     0   | (3221...)|     1        -> unsigned 이므로 0이 출력됨.
        rom[13] = 32'b000000001111_00010_100_01001_0010011;  // xori x9, x2, 15          => 3(0011) | 12(1100) |    15(1111)  
        rom[14] = 32'b000000001111_00010_110_01010_0010011;  // ori  x10, x2, 15         => 15(1111)| 12(1100) |    15(1111)  
        rom[15] = 32'b000000001111_00010_111_01011_0010011;  // andi x11, x2, 15         => 12(1100)| 12(1100) |    15(1111)  

        //rom[x]=32'b funct7 _shamt_ rs1 _f3 _ rd  _ op        // I-TYPE shift (7-bit imm)           rd
        rom[16] = 32'b0000000_10111_00101_001_01100_0010011;   // slli x12, x5, 23            =>  000000000..000
        rom[17] = 32'b0000000_10111_00101_101_01101_0010011;   // srli x13, x5, 23           =>   00..001100....00
        rom[18] = 32'b0000000_01111_00101_101_01110_0010011;   // srli x14, x5, 15           =>   00..001100....00
        rom[19] = 32'b0100000_10111_00101_101_01111_0010011;   // srai x15, x5, 23             => 11111100....00
        // 추후의 값을 합성하기 위한 add 한번 => 위의 rom[17]과 rom[18]을 더하여 값을 생성.
        rom[20] = 32'b0000000_01110_01101_000_10100_0110011;   // add  x20, x13, x14        => 16,17 번쨰와 8,9 번 째 bit가 1인 값 생성.
                                                                                                // 00000000000000011000000110000000

        //rom[x]=32'b  imm7 _ rs2  _ rs1 _ f3_ imm5 _ op       // S-TYPE (store)     주소 계산                    ram_addr   |     rd
        rom[21] = 32'b0000000_10100_00010_000_01000_0100011;  // sb  x20, 8(x2)   -> 12+8=20(5)           =>         5      |   00...00000000000100...0
        rom[22] = 32'b0000000_10100_00010_001_01100_0100011;  // sh  x20, 12(x2)  -> 12+12=24(6)          =>         6      |   00...00010000001100...0
        rom[23] = 32'b0000000_10100_00010_010_10000_0100011;  // sw  x20, 16(x2)  -> 12+16=28(7)          =>         7      |   00...00110000001100...0

        //rom[x]=32'b  imm12      _ rs1 _ f3_ rd  _   op      // L-TYPE (load)      주소 계산       ram_addr     |      rd
        rom[24] = 32'b000000011100_00000_100_01111_0000011;   // lbu  x15, 28(x0)   0+28=28  =>     7           |   00............00   
        rom[25] = 32'b000000011100_00000_000_10000_0000011;   // lb   x16, 28(x0)   0+28=28  =>     7           |   00............00
        rom[26] = 32'b000000011100_00000_101_10001_0000011;   // lhu  x17, 28(x0)   0+28=28  =>     7           |   00...0011000..00             
        rom[27] = 32'b000000011100_00000_001_10010_0000011;   // lh   x18, 28(x0)   0+28=28  =>     7           |   111...111000..00    
        rom[28] = 32'b000000011100_00000_010_10011_0000011;   // lw   x19, 28(x0)   0+28=28  =>     7           |   111...111000..00

        //rom[x]=32'b   imm7 _ rs2 _ rs1 _f3 _imm5 _ opcode      // B-TYPE
        rom[29] = 32'b0000000_00010_00010_000_01100_1100011;      // beq  x2, x2, 12    -> 증가O
        rom[32] = 32'b0000000_00010_00000_001_01100_1100011;      // bnq  x0, x2, 12    -> 증가O
        rom[35] = 32'b0000000_00000_00101_100_01100_1100011;      // blt  x5, x0, 12    -> 이 떄는 증가O -> x5를 signed로 읽으면 음수가 되므로.
        rom[38] = 32'b0000000_00000_00101_101_01100_1100011;      // bge  x5, x0, 12    -> 이 때는 증가X -> (위와 동일한 이유)  
        rom[39] = 32'b0000000_00000_00101_110_01100_1100011;      // bltu x5, x0, 12   -> 이 때는 증가X
        rom[40] = 32'b0000000_00000_00101_111_01100_1100011;      // bgeu x5, x0, 12   -> 이 때는 증가O

        //rom[x]= 32'b        imm20       _ rd  _ op        // Upper(LUI & AUIPC)          
        rom[43] = 32'b00000000000000000011_01010_0110111;   // lui   x10, 3  (check!) ->  0000000000000000_0011000000000000 가 RF에 저장됨.
        rom[44] = 32'b00000000000000000000_01011_0010111;   // auipc x11, 0  (check!) ->  PC : 44 * 4 = 176 -> rd에 176이 저장되도록 함!
        
        // jal에서는 imm의 배열 순서가 뒤죽박죽인 것에 주의.
        //  imm[20][10:1][11][19:12]
        // imm[0]=0은 별도로 DataPath에서 설정         
        //rom[x]= 32'b      imm(20)       _ rd  _ op        // Jump And Link
        rom[45] = 32'b00000000110000000000_01100_1101111;   // jal   x12, 12           ->  PC = 45 * 4 = 180 -> rd = PC + 4 = 184, PC = PC + imm = 180 + 12 = 192
        
        //rom[x]= 32'b   imm(12)  _ rs1 _f3 _ rd  _  op
        rom[48] = 32'b000000010000_01100_000_01101_1100111; // jalr x13, x12, 16        -> PC = 48 * 4 = 192 -> rd = PC + 4 = 196, PC = rs1 + imm = 184 + 16 = 200
    end               

    assign data = rom[addr[31:2]];
 
endmodule



